module mod_a ( input in1, input in2, output out );
    // Module body
    // Since this is an example we will use and OR gate 
    assign out = in1 | in2;

endmodule